`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:26:30 05/07/2018 
// Design Name: 
// Module Name:    sim_test_girovettori 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module sim_test_girovettori(
		input [10:0] in,
		output reg [0:10] out
    );

assign out = 11'd6;

endmodule
